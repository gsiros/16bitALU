library verilog;
use verilog.vl_types.all;
entity ErgasiaDyo_vlg_vec_tst is
end ErgasiaDyo_vlg_vec_tst;
